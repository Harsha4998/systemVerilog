module test_event;
  logic addr;
  logic data;
  initial begin 
  end
endmodule
